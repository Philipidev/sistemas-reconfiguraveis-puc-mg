library IEEE;
use IEEE.STD_LOGIC_1164.ALL;  -- Biblioteca para uso de tipos l�gicos padr�o
use IEEE.NUMERIC_STD.ALL;  -- Biblioteca para convers�es num�ricas e opera��es com std_logic_vector

entity RegBank is
    Port (
        clk_in        : in  std_logic;
        nrst          : in  std_logic;
        regn_di       : in  std_logic_vector(7 downto 0);
        regn_wr_sel   : in  std_logic_vector(2 downto 0);
        regn_wr_ena   : in  std_logic;
        regn_rd_sel_a : in  std_logic_vector(2 downto 0);
        regn_rd_sel_b : in  std_logic_vector(2 downto 0);
        c_flag_in     : in  std_logic;
        z_flag_in     : in  std_logic;
        v_flag_in     : in  std_logic;
        c_flag_wr_ena : in  std_logic;
        z_flag_wr_ena : in  std_logic;
        v_flag_wr_ena : in  std_logic;
        regn_do_a     : out std_logic_vector(7 downto 0);
        regn_do_b     : out std_logic_vector(7 downto 0);
        c_flag_out    : out std_logic;
        z_flag_out    : out std_logic;
        v_flag_out    : out std_logic
    );
end RegBank;

architecture Behavioral of RegBank is
    type reg_array is array (7 downto 0) of std_logic_vector(7 downto 0);
    signal regs : reg_array := (others => (others => '0'));
    signal c_flag, z_flag, v_flag : std_logic := '0';
begin
    process(clk_in, nrst)
    begin
        if nrst = '0' then
            regs <= (others => (others => '0'));
            c_flag <= '0';
            z_flag <= '0';
            v_flag <= '0';
        elsif rising_edge(clk_in) then
            -- Write to general registers
            if regn_wr_ena = '1' then
                regs(to_integer(unsigned(regn_wr_sel))) <= regn_di;
            end if;

            -- Write to flags with priority
            if c_flag_wr_ena = '1' then
                regs(7)(0) <= c_flag_in;
            end if;
            if z_flag_wr_ena = '1' then
                regs(7)(1) <= z_flag_in;
            end if;
            if v_flag_wr_ena = '1' then
                regs(7)(2) <= v_flag_in;
            end if;
        end if;
    end process;

    -- Asynchronous read
    regn_do_a <= regs(to_integer(unsigned(regn_rd_sel_a)));
    regn_do_b <= regs(to_integer(unsigned(regn_rd_sel_b)));

    -- Outputs for flags
    c_flag_out <= regs(7)(0);
    z_flag_out <= regs(7)(1);
    v_flag_out <= regs(7)(2);
end Behavioral;
